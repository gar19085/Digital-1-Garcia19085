//Universidad del Valle de Guatemala
//Lab08
//ALU de 4 bits
//Gar19085

module  ALU(A, B, SEL, OUT);
    input   [3:0] A, B;
    input   [:] ;
    output  OUT;  


    case ()
        : 
        default: 
    endcase

endmodule    




