

module testbench();

reg ;
wire ;


ROM4Kx8 Ju87();

initial begin
        $display("\n");
        $display("Ejercicio 2");
        $display("CLK");
        $monitor("%b", CLK);
end


endmodule