//UNIVERSIDAD DEL VALLE 
//LAB09
//Rodrigo GArcía19085


module  ROM4Kx8(address, Dout);
    input   [11:0] address;
    output  [7:0] Dout;

endmodule    