//testbench



module  testbench();



enmodule    