//Universidad del Valle de Guatemala
//Digital 1
//Laboratorio 05
//Rodrigo José García Ambrosy. Carnet: 19085

//Implemento mmódulo Mux 2:1 
module Mux2x1(input wire A, B, SEL, Gbar, output wire Y);
//ands
wire a1, a2;
//nots
wire n1;

//operadores del mux2:1
not(n1, );
and(a1, );
and(a2, );
or(Y, );